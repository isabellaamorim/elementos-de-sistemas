-- Elementos de Sistemas
-- developed by Luciano Soares
-- tb_Ram8.vhd
-- date: 4/4/2017

Library ieee;
use ieee.std_logic_1164.all;

library vunit_lib;
context vunit_lib.vunit_context;

entity tb_Ram8 is
  generic (runner_cfg : string);
end entity;

architecture tb of tb_Ram8 is

	component  Ram8 is
		port(
			clock:   in  STD_LOGIC;
			input:   in  STD_LOGIC_VECTOR(15 downto 0);
			load:    in  STD_LOGIC;
			address: in  STD_LOGIC_VECTOR( 2 downto 0);
			output:  out STD_LOGIC_VECTOR(15 downto 0)
		);
	end component;

	signal inClock : std_logic := '0';
	signal inInput : STD_LOGIC_VECTOR(15 downto 0);
	signal inLoad : STD_LOGIC;
	signal inAddress : STD_LOGIC_VECTOR( 2 downto 0);
	signal outOutput : STD_LOGIC_VECTOR(15 downto 0);

begin

	mapping: Ram8 port map(inClock, inInput, inLoad, inAddress, outOutput);

	inClock <= not inClock after 100 ps;

  main : process
  begin
    test_runner_setup(runner, runner_cfg);

		-- Teste: 0
		inInput <= x"5555"; inAddress <= "000"; inLoad <= '1';
    wait until inClock'event and inClock='0';
		assert(outOutput = x"5555")  report "Falha em teste: 0" severity error;

		-- Teste: 1
		inInput <= x"AAAA"; inAddress <= "000"; inLoad <= '0';
    wait until inClock'event and inClock='0';
		assert(outOutput = x"5555")  report "Falha em teste: 1" severity error;

    -- Teste: 2
		inInput <= x"AAAA"; inAddress <= "010"; inLoad <= '1';
    wait until inClock'event and inClock='0';
		assert(outOutput = x"AAAA")  report "Falha em teste: 1" severity error;

    -- Teste: 3
		inInput <= x"FFFF"; inAddress <= "010"; inLoad <= '0';
    wait until inClock'event and inClock='0';
		assert(outOutput = x"AAAA")  report "Falha em teste: 1" severity error;

    -- Teste: 4
		inInput <= x"FFFF"; inAddress <= "111"; inLoad <= '1';
    wait until inClock'event and inClock='0';
		assert(outOutput = x"FFFF")  report "Falha em teste: 1" severity error;

    -- Teste: 5
		inInput <= x"F0F0"; inAddress <= "111"; inLoad <= '0';
    wait until inClock'event and inClock='0';
		assert(outOutput = x"FFFF")  report "Falha em teste: 1" severity error;

    -- finish
    wait until inClock'event and inClock='0';
    test_runner_cleanup(runner); -- Simulation ends here

	wait;
  end process;
end architecture;
